-- ============================================================================
--   Ver  :| Author            :| Mod. Date :| Changes Made:
--   V1.0 :| T. Rampone        :| 04/09/2017:| -
-- ============================================================================

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.all;

entity DE0_nano_top_level is
	port(	-- CLOCK 50 MHz
			CLOCK_50 :			  in std_logic;
			-- DRAM
			DRAM_ADDR :			  out std_logic_vector(12 downto 0);
			DRAM_BA :			  out std_logic_vector(1 downto 0);
			DRAM_CAS_N :		  out std_logic;
			DRAM_CKE :			  out std_logic;
			DRAM_CLK :			  out std_logic;
			DRAM_CS_N :			  out std_logic;
			DRAM_DQ :			  inout std_logic_vector(15 downto 0);
			DRAM_DQM :			  out std_logic_vector(1 downto 0);
			DRAM_RAS_N :		  out std_logic;
			DRAM_WE_N :			  out std_logic;
			-- KEY
			KEY :				     in std_logic_vector(1 downto 0);
			-- LED
			LED :				     out std_logic_vector(7 downto 0);
         -- SWITCH
			SW :                in std_logic_vector(3 downto 0);
			-- EPCS
			EPCS_DCLK :         out std_logic;
			EPCS_NCSO :         out std_logic;
			EPCS_ASDO :         out std_logic;
			EPCS_DATA0 :        in std_logic;
			-- G SENSOR
			G_SENSOR_CS_N :     out std_logic;
			G_SENSOR_INT :      in std_logic;
			-- EXT SENSOR
			EXT_SENSOR_INT :    in std_logic;
			-- ZigBee
			Xbee_Out :          in std_logic;           -- Xbee_Out -> Rx (to UART)
			Xbee_In :           out std_logic;          -- Xbee_In -> Tx (from UART)
			-- ADC
			ADC_SDAT :          in std_logic;
			ADC_SADDR :         out std_logic;
			ADC_SCLK :          out std_logic;
			ADC_CS_N :          out std_logic;
			-- I2C (internal: DE0-nano)
			I2C_SCLK :          out std_logic;
			I2C_SDAT :          inout std_logic;
			-- I2C (external: extension board with sensors)
			I2C_EXT_SCLK :      out std_logic;
			I2C_EXT_SDA :       inout std_logic;
			-- Arduino interface (digital signals only)
			ARDUINO_IO :        inout std_logic_vector(15 downto 0);
			ARDUINO_RESET_N :   inout std_logic
	);
end DE0_nano_top_level;


architecture rtl of DE0_nano_top_level is
-- pll
signal pll_locked : std_logic;

--I2C
signal i2c_clk : std_logic;

-- System module QSys
component DE0_nano_system is
        port (
            altpll_sys_c1_clk                : out   std_logic;                                        -- clk
            altpll_sys_locked_conduit_export : out   std_logic;                                        -- export
            clk_clk                          : in    std_logic                     := 'X';             -- clk
            epcs_dclk                        : out   std_logic;                                        -- dclk
            epcs_sce                         : out   std_logic;                                        -- sce
            epcs_sdo                         : out   std_logic;                                        -- sdo
            epcs_data0                       : in    std_logic                     := 'X';             -- data0
            g_sensor_irq_export              : in    std_logic                     := 'X';             -- export
            i2c_ext_sda_export               : inout std_logic                     := 'X';             -- export
            i2c_scl_export                   : out   std_logic;                                        -- export
            i2c_sda_export                   : inout std_logic                     := 'X';             -- export
            ext_sensor_irq_export            : in    std_logic                     := 'X';             -- export
            pio_key_export                   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- export
            pio_leds_export                  : out   std_logic_vector(7 downto 0);                     -- export
            pio_switch_export                : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- export
            sdram_wire_addr                  : out   std_logic_vector(12 downto 0);                    -- addr
            sdram_wire_ba                    : out   std_logic_vector(1 downto 0);                     -- ba
            sdram_wire_cas_n                 : out   std_logic;                                        -- cas_n
            sdram_wire_cke                   : out   std_logic;                                        -- cke
            sdram_wire_cs_n                  : out   std_logic;                                        -- cs_n
            sdram_wire_dq                    : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
            sdram_wire_dqm                   : out   std_logic_vector(1 downto 0);                     -- dqm
            sdram_wire_ras_n                 : out   std_logic;                                        -- ras_n
            sdram_wire_we_n                  : out   std_logic;                                        -- we_n
            reset_reset_n                    : in    std_logic;                                        -- reset_n
            xbee_rxd                      	: in    std_logic                     := 'X';             -- rxd
            xbee_txd                      	: out   std_logic;                                        -- txd
            adc_spi_conduit_MISO             : in    std_logic                     := 'X';             -- MISO
            adc_spi_conduit_MOSI             : out   std_logic;                                        -- MOSI
            adc_spi_conduit_SCLK             : out   std_logic;                                        -- SCLK
            adc_spi_conduit_SS_n             : out   std_logic                                         -- SS_n
            );
end component DE0_nano_system;

begin
-- G SENSOR
G_SENSOR_CS_N <= '1';

-- I2C clk
I2C_SCLK <= i2c_clk;
I2C_EXT_SCLK <= i2c_clk;

-- QSys module 
u0 : component DE0_nano_system
    port map (
            altpll_sys_c1_clk                => DRAM_CLK,
            altpll_sys_locked_conduit_export => pll_locked,
            clk_clk                          => CLOCK_50,
            epcs_dclk                        => EPCS_DCLK,
            epcs_sce                         => EPCS_NCSO,
            epcs_sdo                         => EPCS_ASDO,
            epcs_data0                       => EPCS_DATA0,
            g_sensor_irq_export              => G_SENSOR_INT,
            i2c_ext_sda_export               => I2C_EXT_SDA,
            i2c_scl_export                   => i2c_clk,            --common to internal and external i2c bus
            i2c_sda_export                   => I2C_SDAT,
            ext_sensor_irq_export            => EXT_SENSOR_INT,
            pio_key_export                   => KEY,
            pio_leds_export                  => LED,
            pio_switch_export                => SW,
            sdram_wire_addr                  => DRAM_ADDR,
            sdram_wire_ba                    => DRAM_BA,
            sdram_wire_cas_n                 => DRAM_CAS_N,
            sdram_wire_cke                   => DRAM_CKE,
            sdram_wire_cs_n                  => DRAM_CS_N,
            sdram_wire_dq                    => DRAM_DQ,
            sdram_wire_dqm                   => DRAM_DQM,
            sdram_wire_ras_n                 => DRAM_RAS_N,
            sdram_wire_we_n                  => DRAM_WE_N,
            reset_reset_n                    => ARDUINO_RESET_N,                 --                          .we_n
            xbee_rxd                      	=> Xbee_Out,                      	--                   tx_xbee.rxd
            xbee_txd                      	=> Xbee_In,                      	--                          .txd
            adc_spi_conduit_MISO             => ADC_SDAT,             				--           adc_spi_conduit.MISO
            adc_spi_conduit_MOSI             => ADC_SADDR,             				--                          .MOSI
            adc_spi_conduit_SCLK             => ADC_SCLK,             				--                          .SCLK
            adc_spi_conduit_SS_n             => ADC_CS_N     
    );

end architecture rtl;