-- DE0_nano_system.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DE0_nano_system is
	port (
		adc_spi_conduit_MISO             : in    std_logic                     := '0';             --           adc_spi_conduit.MISO
		adc_spi_conduit_MOSI             : out   std_logic;                                        --                          .MOSI
		adc_spi_conduit_SCLK             : out   std_logic;                                        --                          .SCLK
		adc_spi_conduit_SS_n             : out   std_logic;                                        --                          .SS_n
		altpll_sys_c1_clk                : out   std_logic;                                        --             altpll_sys_c1.clk
		altpll_sys_locked_conduit_export : out   std_logic;                                        -- altpll_sys_locked_conduit.export
		clk_clk                          : in    std_logic                     := '0';             --                       clk.clk
		epcs_dclk                        : out   std_logic;                                        --                      epcs.dclk
		epcs_sce                         : out   std_logic;                                        --                          .sce
		epcs_sdo                         : out   std_logic;                                        --                          .sdo
		epcs_data0                       : in    std_logic                     := '0';             --                          .data0
		ext_sensor_irq_export            : in    std_logic                     := '0';             --            ext_sensor_irq.export
		g_sensor_irq_export              : in    std_logic                     := '0';             --              g_sensor_irq.export
		i2c_ext_sda_export               : inout std_logic                     := '0';             --               i2c_ext_sda.export
		i2c_scl_export                   : out   std_logic;                                        --                   i2c_scl.export
		i2c_sda_export                   : inout std_logic                     := '0';             --                   i2c_sda.export
		pio_key_export                   : in    std_logic_vector(1 downto 0)  := (others => '0'); --                   pio_key.export
		pio_leds_export                  : out   std_logic_vector(7 downto 0);                     --                  pio_leds.export
		pio_switch_export                : in    std_logic_vector(3 downto 0)  := (others => '0'); --                pio_switch.export
		reset_reset_n                    : in    std_logic                     := '0';             --                     reset.reset_n
		sdram_wire_addr                  : out   std_logic_vector(12 downto 0);                    --                sdram_wire.addr
		sdram_wire_ba                    : out   std_logic_vector(1 downto 0);                     --                          .ba
		sdram_wire_cas_n                 : out   std_logic;                                        --                          .cas_n
		sdram_wire_cke                   : out   std_logic;                                        --                          .cke
		sdram_wire_cs_n                  : out   std_logic;                                        --                          .cs_n
		sdram_wire_dq                    : inout std_logic_vector(15 downto 0) := (others => '0'); --                          .dq
		sdram_wire_dqm                   : out   std_logic_vector(1 downto 0);                     --                          .dqm
		sdram_wire_ras_n                 : out   std_logic;                                        --                          .ras_n
		sdram_wire_we_n                  : out   std_logic;                                        --                          .we_n
		xbee_rxd                         : in    std_logic                     := '0';             --                      xbee.rxd
		xbee_txd                         : out   std_logic                                         --                          .txd
	);
end entity DE0_nano_system;

architecture rtl of DE0_nano_system is
	component DE0_nano_system_adc_spi_int is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component DE0_nano_system_adc_spi_int;

	component DE0_nano_system_altpll_sys is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			locked             : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X';             -- export
			areset             : in  std_logic                     := 'X';             -- export
			phasedone          : out std_logic                                         -- export
		);
	end component DE0_nano_system_altpll_sys;

	component altera_avalon_mm_clock_crossing_bridge is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			HDL_ADDR_WIDTH      : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             -- clk
			m0_reset         : in  std_logic                     := 'X';             -- reset
			s0_clk           : in  std_logic                     := 'X';             -- clk
			s0_reset         : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(11 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component altera_avalon_mm_clock_crossing_bridge;

	component DE0_nano_system_epcs is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			address    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read_n     : in  std_logic                     := 'X';             -- read_n
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			irq        : out std_logic;                                        -- irq
			dclk       : out std_logic;                                        -- export
			sce        : out std_logic;                                        -- export
			sdo        : out std_logic;                                        -- export
			data0      : in  std_logic                     := 'X'              -- export
		);
	end component DE0_nano_system_epcs;

	component DE0_nano_system_ext_sensor_int is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component DE0_nano_system_ext_sensor_int;

	component DE0_nano_system_g_sensor_int is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component DE0_nano_system_g_sensor_int;

	component DE0_nano_system_i2c_EXT_sda is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic                     := 'X'              -- export
		);
	end component DE0_nano_system_i2c_EXT_sda;

	component DE0_nano_system_i2c_scl is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component DE0_nano_system_i2c_scl;

	component DE0_nano_system_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component DE0_nano_system_jtag_uart;

	component DE0_nano_system_nios2_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component DE0_nano_system_nios2_cpu;

	component DE0_nano_system_onchip_mem is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component DE0_nano_system_onchip_mem;

	component DE0_nano_system_pio_key is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component DE0_nano_system_pio_key;

	component DE0_nano_system_pio_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component DE0_nano_system_pio_leds;

	component DE0_nano_system_pio_switch is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component DE0_nano_system_pio_switch;

	component DE0_nano_system_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component DE0_nano_system_sdram;

	component DE0_nano_system_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component DE0_nano_system_sysid_qsys;

	component DE0_nano_system_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component DE0_nano_system_timer;

	component DE0_nano_system_xbee_uart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component DE0_nano_system_xbee_uart;

	component DE0_nano_system_mm_interconnect_0 is
		port (
			altpll_sys_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			clk_50_clk_clk                                               : in  std_logic                     := 'X';             -- clk
			altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_cpu_reset_reset_bridge_in_reset_reset                  : in  std_logic                     := 'X';             -- reset
			nios2_cpu_data_master_address                                : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_cpu_data_master_waitrequest                            : out std_logic;                                        -- waitrequest
			nios2_cpu_data_master_byteenable                             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_cpu_data_master_read                                   : in  std_logic                     := 'X';             -- read
			nios2_cpu_data_master_readdata                               : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_cpu_data_master_readdatavalid                          : out std_logic;                                        -- readdatavalid
			nios2_cpu_data_master_write                                  : in  std_logic                     := 'X';             -- write
			nios2_cpu_data_master_writedata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_cpu_data_master_debugaccess                            : in  std_logic                     := 'X';             -- debugaccess
			nios2_cpu_instruction_master_address                         : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_cpu_instruction_master_waitrequest                     : out std_logic;                                        -- waitrequest
			nios2_cpu_instruction_master_read                            : in  std_logic                     := 'X';             -- read
			nios2_cpu_instruction_master_readdata                        : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_cpu_instruction_master_readdatavalid                   : out std_logic;                                        -- readdatavalid
			altpll_sys_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			altpll_sys_pll_slave_write                                   : out std_logic;                                        -- write
			altpll_sys_pll_slave_read                                    : out std_logic;                                        -- read
			altpll_sys_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_sys_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			clock_crossing_bridge_IO_s0_address                          : out std_logic_vector(11 downto 0);                    -- address
			clock_crossing_bridge_IO_s0_write                            : out std_logic;                                        -- write
			clock_crossing_bridge_IO_s0_read                             : out std_logic;                                        -- read
			clock_crossing_bridge_IO_s0_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			clock_crossing_bridge_IO_s0_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			clock_crossing_bridge_IO_s0_burstcount                       : out std_logic_vector(0 downto 0);                     -- burstcount
			clock_crossing_bridge_IO_s0_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			clock_crossing_bridge_IO_s0_readdatavalid                    : in  std_logic                     := 'X';             -- readdatavalid
			clock_crossing_bridge_IO_s0_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			clock_crossing_bridge_IO_s0_debugaccess                      : out std_logic;                                        -- debugaccess
			jtag_uart_avalon_jtag_slave_address                          : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                            : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                             : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                       : out std_logic;                                        -- chipselect
			nios2_cpu_debug_mem_slave_address                            : out std_logic_vector(8 downto 0);                     -- address
			nios2_cpu_debug_mem_slave_write                              : out std_logic;                                        -- write
			nios2_cpu_debug_mem_slave_read                               : out std_logic;                                        -- read
			nios2_cpu_debug_mem_slave_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_cpu_debug_mem_slave_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_cpu_debug_mem_slave_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_cpu_debug_mem_slave_waitrequest                        : in  std_logic                     := 'X';             -- waitrequest
			nios2_cpu_debug_mem_slave_debugaccess                        : out std_logic;                                        -- debugaccess
			onchip_mem_s1_address                                        : out std_logic_vector(9 downto 0);                     -- address
			onchip_mem_s1_write                                          : out std_logic;                                        -- write
			onchip_mem_s1_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_mem_s1_writedata                                      : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_mem_s1_byteenable                                     : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_mem_s1_chipselect                                     : out std_logic;                                        -- chipselect
			onchip_mem_s1_clken                                          : out std_logic;                                        -- clken
			sdram_s1_address                                             : out std_logic_vector(23 downto 0);                    -- address
			sdram_s1_write                                               : out std_logic;                                        -- write
			sdram_s1_read                                                : out std_logic;                                        -- read
			sdram_s1_readdata                                            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                                           : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                                          : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                                       : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                                         : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                                          : out std_logic                                         -- chipselect
		);
	end component DE0_nano_system_mm_interconnect_0;

	component DE0_nano_system_mm_interconnect_1 is
		port (
			altpll_sys_c2_clk                                             : in  std_logic                     := 'X';             -- clk
			clock_crossing_bridge_IO_m0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			clock_crossing_bridge_IO_m0_address                           : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clock_crossing_bridge_IO_m0_waitrequest                       : out std_logic;                                        -- waitrequest
			clock_crossing_bridge_IO_m0_burstcount                        : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			clock_crossing_bridge_IO_m0_byteenable                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clock_crossing_bridge_IO_m0_read                              : in  std_logic                     := 'X';             -- read
			clock_crossing_bridge_IO_m0_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			clock_crossing_bridge_IO_m0_readdatavalid                     : out std_logic;                                        -- readdatavalid
			clock_crossing_bridge_IO_m0_write                             : in  std_logic                     := 'X';             -- write
			clock_crossing_bridge_IO_m0_writedata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			clock_crossing_bridge_IO_m0_debugaccess                       : in  std_logic                     := 'X';             -- debugaccess
			adc_spi_int_spi_control_port_address                          : out std_logic_vector(2 downto 0);                     -- address
			adc_spi_int_spi_control_port_write                            : out std_logic;                                        -- write
			adc_spi_int_spi_control_port_read                             : out std_logic;                                        -- read
			adc_spi_int_spi_control_port_readdata                         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			adc_spi_int_spi_control_port_writedata                        : out std_logic_vector(15 downto 0);                    -- writedata
			adc_spi_int_spi_control_port_chipselect                       : out std_logic;                                        -- chipselect
			epcs_epcs_control_port_address                                : out std_logic_vector(8 downto 0);                     -- address
			epcs_epcs_control_port_write                                  : out std_logic;                                        -- write
			epcs_epcs_control_port_read                                   : out std_logic;                                        -- read
			epcs_epcs_control_port_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			epcs_epcs_control_port_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			epcs_epcs_control_port_chipselect                             : out std_logic;                                        -- chipselect
			ext_sensor_int_s1_address                                     : out std_logic_vector(1 downto 0);                     -- address
			ext_sensor_int_s1_write                                       : out std_logic;                                        -- write
			ext_sensor_int_s1_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ext_sensor_int_s1_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			ext_sensor_int_s1_chipselect                                  : out std_logic;                                        -- chipselect
			g_sensor_int_s1_address                                       : out std_logic_vector(1 downto 0);                     -- address
			g_sensor_int_s1_write                                         : out std_logic;                                        -- write
			g_sensor_int_s1_readdata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			g_sensor_int_s1_writedata                                     : out std_logic_vector(31 downto 0);                    -- writedata
			g_sensor_int_s1_chipselect                                    : out std_logic;                                        -- chipselect
			i2c_EXT_sda_s1_address                                        : out std_logic_vector(1 downto 0);                     -- address
			i2c_EXT_sda_s1_write                                          : out std_logic;                                        -- write
			i2c_EXT_sda_s1_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i2c_EXT_sda_s1_writedata                                      : out std_logic_vector(31 downto 0);                    -- writedata
			i2c_EXT_sda_s1_chipselect                                     : out std_logic;                                        -- chipselect
			i2c_scl_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			i2c_scl_s1_write                                              : out std_logic;                                        -- write
			i2c_scl_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i2c_scl_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			i2c_scl_s1_chipselect                                         : out std_logic;                                        -- chipselect
			i2c_sda_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			i2c_sda_s1_write                                              : out std_logic;                                        -- write
			i2c_sda_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i2c_sda_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			i2c_sda_s1_chipselect                                         : out std_logic;                                        -- chipselect
			pio_key_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			pio_key_s1_write                                              : out std_logic;                                        -- write
			pio_key_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_key_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			pio_key_s1_chipselect                                         : out std_logic;                                        -- chipselect
			pio_leds_s1_address                                           : out std_logic_vector(1 downto 0);                     -- address
			pio_leds_s1_write                                             : out std_logic;                                        -- write
			pio_leds_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_leds_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			pio_leds_s1_chipselect                                        : out std_logic;                                        -- chipselect
			pio_switch_s1_address                                         : out std_logic_vector(1 downto 0);                     -- address
			pio_switch_s1_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sysid_qsys_control_slave_address                              : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_control_slave_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_s1_address                                              : out std_logic_vector(2 downto 0);                     -- address
			timer_s1_write                                                : out std_logic;                                        -- write
			timer_s1_readdata                                             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_s1_writedata                                            : out std_logic_vector(15 downto 0);                    -- writedata
			timer_s1_chipselect                                           : out std_logic;                                        -- chipselect
			xbee_uart_s1_address                                          : out std_logic_vector(2 downto 0);                     -- address
			xbee_uart_s1_write                                            : out std_logic;                                        -- write
			xbee_uart_s1_read                                             : out std_logic;                                        -- read
			xbee_uart_s1_readdata                                         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			xbee_uart_s1_writedata                                        : out std_logic_vector(15 downto 0);                    -- writedata
			xbee_uart_s1_begintransfer                                    : out std_logic;                                        -- begintransfer
			xbee_uart_s1_chipselect                                       : out std_logic                                         -- chipselect
		);
	end component DE0_nano_system_mm_interconnect_1;

	component DE0_nano_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			receiver6_irq : in  std_logic                     := 'X'; -- irq
			receiver7_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component DE0_nano_system_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component de0_nano_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component de0_nano_system_rst_controller;

	component de0_nano_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component de0_nano_system_rst_controller_001;

	signal altpll_sys_c0_clk                                              : std_logic;                     -- altpll_sys:c0 -> [clock_crossing_bridge_IO:s0_clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, irq_synchronizer_004:sender_clk, irq_synchronizer_005:sender_clk, irq_synchronizer_006:sender_clk, jtag_uart:clk, mm_interconnect_0:altpll_sys_c0_clk, nios2_cpu:clk, onchip_mem:clk, rst_controller_002:clk, sdram:clk]
	signal altpll_sys_c2_clk                                              : std_logic;                     -- altpll_sys:c2 -> [adc_spi_int:clk, clock_crossing_bridge_IO:m0_clk, epcs:clk, ext_sensor_int:clk, g_sensor_int:clk, i2c_EXT_sda:clk, i2c_scl:clk, i2c_sda:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, irq_synchronizer_003:receiver_clk, irq_synchronizer_004:receiver_clk, irq_synchronizer_005:receiver_clk, irq_synchronizer_006:receiver_clk, mm_interconnect_1:altpll_sys_c2_clk, pio_key:clk, pio_leds:clk, pio_switch:clk, rst_controller:clk, sysid_qsys:clock, timer:clk, xbee_uart:clk]
	signal nios2_cpu_data_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_cpu_data_master_readdata -> nios2_cpu:d_readdata
	signal nios2_cpu_data_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:nios2_cpu_data_master_waitrequest -> nios2_cpu:d_waitrequest
	signal nios2_cpu_data_master_debugaccess                              : std_logic;                     -- nios2_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_cpu_data_master_debugaccess
	signal nios2_cpu_data_master_address                                  : std_logic_vector(26 downto 0); -- nios2_cpu:d_address -> mm_interconnect_0:nios2_cpu_data_master_address
	signal nios2_cpu_data_master_byteenable                               : std_logic_vector(3 downto 0);  -- nios2_cpu:d_byteenable -> mm_interconnect_0:nios2_cpu_data_master_byteenable
	signal nios2_cpu_data_master_read                                     : std_logic;                     -- nios2_cpu:d_read -> mm_interconnect_0:nios2_cpu_data_master_read
	signal nios2_cpu_data_master_readdatavalid                            : std_logic;                     -- mm_interconnect_0:nios2_cpu_data_master_readdatavalid -> nios2_cpu:d_readdatavalid
	signal nios2_cpu_data_master_write                                    : std_logic;                     -- nios2_cpu:d_write -> mm_interconnect_0:nios2_cpu_data_master_write
	signal nios2_cpu_data_master_writedata                                : std_logic_vector(31 downto 0); -- nios2_cpu:d_writedata -> mm_interconnect_0:nios2_cpu_data_master_writedata
	signal nios2_cpu_instruction_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_cpu_instruction_master_readdata -> nios2_cpu:i_readdata
	signal nios2_cpu_instruction_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:nios2_cpu_instruction_master_waitrequest -> nios2_cpu:i_waitrequest
	signal nios2_cpu_instruction_master_address                           : std_logic_vector(26 downto 0); -- nios2_cpu:i_address -> mm_interconnect_0:nios2_cpu_instruction_master_address
	signal nios2_cpu_instruction_master_read                              : std_logic;                     -- nios2_cpu:i_read -> mm_interconnect_0:nios2_cpu_instruction_master_read
	signal nios2_cpu_instruction_master_readdatavalid                     : std_logic;                     -- mm_interconnect_0:nios2_cpu_instruction_master_readdatavalid -> nios2_cpu:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect       : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata         : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest      : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address          : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read             : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata           : std_logic_vector(31 downto 0); -- nios2_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios2_cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest        : std_logic;                     -- nios2_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess        : std_logic;                     -- mm_interconnect_0:nios2_cpu_debug_mem_slave_debugaccess -> nios2_cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_address            : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_cpu_debug_mem_slave_address -> nios2_cpu:debug_mem_slave_address
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_read               : std_logic;                     -- mm_interconnect_0:nios2_cpu_debug_mem_slave_read -> nios2_cpu:debug_mem_slave_read
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_cpu_debug_mem_slave_byteenable -> nios2_cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_write              : std_logic;                     -- mm_interconnect_0:nios2_cpu_debug_mem_slave_write -> nios2_cpu:debug_mem_slave_write
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_cpu_debug_mem_slave_writedata -> nios2_cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_altpll_sys_pll_slave_readdata                : std_logic_vector(31 downto 0); -- altpll_sys:readdata -> mm_interconnect_0:altpll_sys_pll_slave_readdata
	signal mm_interconnect_0_altpll_sys_pll_slave_address                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:altpll_sys_pll_slave_address -> altpll_sys:address
	signal mm_interconnect_0_altpll_sys_pll_slave_read                    : std_logic;                     -- mm_interconnect_0:altpll_sys_pll_slave_read -> altpll_sys:read
	signal mm_interconnect_0_altpll_sys_pll_slave_write                   : std_logic;                     -- mm_interconnect_0:altpll_sys_pll_slave_write -> altpll_sys:write
	signal mm_interconnect_0_altpll_sys_pll_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:altpll_sys_pll_slave_writedata -> altpll_sys:writedata
	signal mm_interconnect_0_clock_crossing_bridge_io_s0_readdata         : std_logic_vector(31 downto 0); -- clock_crossing_bridge_IO:s0_readdata -> mm_interconnect_0:clock_crossing_bridge_IO_s0_readdata
	signal mm_interconnect_0_clock_crossing_bridge_io_s0_waitrequest      : std_logic;                     -- clock_crossing_bridge_IO:s0_waitrequest -> mm_interconnect_0:clock_crossing_bridge_IO_s0_waitrequest
	signal mm_interconnect_0_clock_crossing_bridge_io_s0_debugaccess      : std_logic;                     -- mm_interconnect_0:clock_crossing_bridge_IO_s0_debugaccess -> clock_crossing_bridge_IO:s0_debugaccess
	signal mm_interconnect_0_clock_crossing_bridge_io_s0_address          : std_logic_vector(11 downto 0); -- mm_interconnect_0:clock_crossing_bridge_IO_s0_address -> clock_crossing_bridge_IO:s0_address
	signal mm_interconnect_0_clock_crossing_bridge_io_s0_read             : std_logic;                     -- mm_interconnect_0:clock_crossing_bridge_IO_s0_read -> clock_crossing_bridge_IO:s0_read
	signal mm_interconnect_0_clock_crossing_bridge_io_s0_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:clock_crossing_bridge_IO_s0_byteenable -> clock_crossing_bridge_IO:s0_byteenable
	signal mm_interconnect_0_clock_crossing_bridge_io_s0_readdatavalid    : std_logic;                     -- clock_crossing_bridge_IO:s0_readdatavalid -> mm_interconnect_0:clock_crossing_bridge_IO_s0_readdatavalid
	signal mm_interconnect_0_clock_crossing_bridge_io_s0_write            : std_logic;                     -- mm_interconnect_0:clock_crossing_bridge_IO_s0_write -> clock_crossing_bridge_IO:s0_write
	signal mm_interconnect_0_clock_crossing_bridge_io_s0_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:clock_crossing_bridge_IO_s0_writedata -> clock_crossing_bridge_IO:s0_writedata
	signal mm_interconnect_0_clock_crossing_bridge_io_s0_burstcount       : std_logic_vector(0 downto 0);  -- mm_interconnect_0:clock_crossing_bridge_IO_s0_burstcount -> clock_crossing_bridge_IO:s0_burstcount
	signal mm_interconnect_0_onchip_mem_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_chipselect -> onchip_mem:chipselect
	signal mm_interconnect_0_onchip_mem_s1_readdata                       : std_logic_vector(31 downto 0); -- onchip_mem:readdata -> mm_interconnect_0:onchip_mem_s1_readdata
	signal mm_interconnect_0_onchip_mem_s1_address                        : std_logic_vector(9 downto 0);  -- mm_interconnect_0:onchip_mem_s1_address -> onchip_mem:address
	signal mm_interconnect_0_onchip_mem_s1_byteenable                     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_mem_s1_byteenable -> onchip_mem:byteenable
	signal mm_interconnect_0_onchip_mem_s1_write                          : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_write -> onchip_mem:write
	signal mm_interconnect_0_onchip_mem_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_mem_s1_writedata -> onchip_mem:writedata
	signal mm_interconnect_0_onchip_mem_s1_clken                          : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_clken -> onchip_mem:clken
	signal mm_interconnect_0_sdram_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                            : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                         : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                             : std_logic_vector(23 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                                : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                       : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                               : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                           : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal clock_crossing_bridge_io_m0_waitrequest                        : std_logic;                     -- mm_interconnect_1:clock_crossing_bridge_IO_m0_waitrequest -> clock_crossing_bridge_IO:m0_waitrequest
	signal clock_crossing_bridge_io_m0_readdata                           : std_logic_vector(31 downto 0); -- mm_interconnect_1:clock_crossing_bridge_IO_m0_readdata -> clock_crossing_bridge_IO:m0_readdata
	signal clock_crossing_bridge_io_m0_debugaccess                        : std_logic;                     -- clock_crossing_bridge_IO:m0_debugaccess -> mm_interconnect_1:clock_crossing_bridge_IO_m0_debugaccess
	signal clock_crossing_bridge_io_m0_address                            : std_logic_vector(11 downto 0); -- clock_crossing_bridge_IO:m0_address -> mm_interconnect_1:clock_crossing_bridge_IO_m0_address
	signal clock_crossing_bridge_io_m0_read                               : std_logic;                     -- clock_crossing_bridge_IO:m0_read -> mm_interconnect_1:clock_crossing_bridge_IO_m0_read
	signal clock_crossing_bridge_io_m0_byteenable                         : std_logic_vector(3 downto 0);  -- clock_crossing_bridge_IO:m0_byteenable -> mm_interconnect_1:clock_crossing_bridge_IO_m0_byteenable
	signal clock_crossing_bridge_io_m0_readdatavalid                      : std_logic;                     -- mm_interconnect_1:clock_crossing_bridge_IO_m0_readdatavalid -> clock_crossing_bridge_IO:m0_readdatavalid
	signal clock_crossing_bridge_io_m0_writedata                          : std_logic_vector(31 downto 0); -- clock_crossing_bridge_IO:m0_writedata -> mm_interconnect_1:clock_crossing_bridge_IO_m0_writedata
	signal clock_crossing_bridge_io_m0_write                              : std_logic;                     -- clock_crossing_bridge_IO:m0_write -> mm_interconnect_1:clock_crossing_bridge_IO_m0_write
	signal clock_crossing_bridge_io_m0_burstcount                         : std_logic_vector(0 downto 0);  -- clock_crossing_bridge_IO:m0_burstcount -> mm_interconnect_1:clock_crossing_bridge_IO_m0_burstcount
	signal mm_interconnect_1_sysid_qsys_control_slave_readdata            : std_logic_vector(31 downto 0); -- sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	signal mm_interconnect_1_sysid_qsys_control_slave_address             : std_logic_vector(0 downto 0);  -- mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	signal mm_interconnect_1_epcs_epcs_control_port_chipselect            : std_logic;                     -- mm_interconnect_1:epcs_epcs_control_port_chipselect -> epcs:chipselect
	signal mm_interconnect_1_epcs_epcs_control_port_readdata              : std_logic_vector(31 downto 0); -- epcs:readdata -> mm_interconnect_1:epcs_epcs_control_port_readdata
	signal mm_interconnect_1_epcs_epcs_control_port_address               : std_logic_vector(8 downto 0);  -- mm_interconnect_1:epcs_epcs_control_port_address -> epcs:address
	signal mm_interconnect_1_epcs_epcs_control_port_read                  : std_logic;                     -- mm_interconnect_1:epcs_epcs_control_port_read -> mm_interconnect_1_epcs_epcs_control_port_read:in
	signal mm_interconnect_1_epcs_epcs_control_port_write                 : std_logic;                     -- mm_interconnect_1:epcs_epcs_control_port_write -> mm_interconnect_1_epcs_epcs_control_port_write:in
	signal mm_interconnect_1_epcs_epcs_control_port_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_1:epcs_epcs_control_port_writedata -> epcs:writedata
	signal mm_interconnect_1_timer_s1_chipselect                          : std_logic;                     -- mm_interconnect_1:timer_s1_chipselect -> timer:chipselect
	signal mm_interconnect_1_timer_s1_readdata                            : std_logic_vector(15 downto 0); -- timer:readdata -> mm_interconnect_1:timer_s1_readdata
	signal mm_interconnect_1_timer_s1_address                             : std_logic_vector(2 downto 0);  -- mm_interconnect_1:timer_s1_address -> timer:address
	signal mm_interconnect_1_timer_s1_write                               : std_logic;                     -- mm_interconnect_1:timer_s1_write -> mm_interconnect_1_timer_s1_write:in
	signal mm_interconnect_1_timer_s1_writedata                           : std_logic_vector(15 downto 0); -- mm_interconnect_1:timer_s1_writedata -> timer:writedata
	signal mm_interconnect_1_pio_leds_s1_chipselect                       : std_logic;                     -- mm_interconnect_1:pio_leds_s1_chipselect -> pio_leds:chipselect
	signal mm_interconnect_1_pio_leds_s1_readdata                         : std_logic_vector(31 downto 0); -- pio_leds:readdata -> mm_interconnect_1:pio_leds_s1_readdata
	signal mm_interconnect_1_pio_leds_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_1:pio_leds_s1_address -> pio_leds:address
	signal mm_interconnect_1_pio_leds_s1_write                            : std_logic;                     -- mm_interconnect_1:pio_leds_s1_write -> mm_interconnect_1_pio_leds_s1_write:in
	signal mm_interconnect_1_pio_leds_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_1:pio_leds_s1_writedata -> pio_leds:writedata
	signal mm_interconnect_1_pio_key_s1_chipselect                        : std_logic;                     -- mm_interconnect_1:pio_key_s1_chipselect -> pio_key:chipselect
	signal mm_interconnect_1_pio_key_s1_readdata                          : std_logic_vector(31 downto 0); -- pio_key:readdata -> mm_interconnect_1:pio_key_s1_readdata
	signal mm_interconnect_1_pio_key_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_1:pio_key_s1_address -> pio_key:address
	signal mm_interconnect_1_pio_key_s1_write                             : std_logic;                     -- mm_interconnect_1:pio_key_s1_write -> mm_interconnect_1_pio_key_s1_write:in
	signal mm_interconnect_1_pio_key_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_1:pio_key_s1_writedata -> pio_key:writedata
	signal mm_interconnect_1_pio_switch_s1_readdata                       : std_logic_vector(31 downto 0); -- pio_switch:readdata -> mm_interconnect_1:pio_switch_s1_readdata
	signal mm_interconnect_1_pio_switch_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_1:pio_switch_s1_address -> pio_switch:address
	signal mm_interconnect_1_g_sensor_int_s1_chipselect                   : std_logic;                     -- mm_interconnect_1:g_sensor_int_s1_chipselect -> g_sensor_int:chipselect
	signal mm_interconnect_1_g_sensor_int_s1_readdata                     : std_logic_vector(31 downto 0); -- g_sensor_int:readdata -> mm_interconnect_1:g_sensor_int_s1_readdata
	signal mm_interconnect_1_g_sensor_int_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_1:g_sensor_int_s1_address -> g_sensor_int:address
	signal mm_interconnect_1_g_sensor_int_s1_write                        : std_logic;                     -- mm_interconnect_1:g_sensor_int_s1_write -> mm_interconnect_1_g_sensor_int_s1_write:in
	signal mm_interconnect_1_g_sensor_int_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_1:g_sensor_int_s1_writedata -> g_sensor_int:writedata
	signal mm_interconnect_1_i2c_sda_s1_chipselect                        : std_logic;                     -- mm_interconnect_1:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	signal mm_interconnect_1_i2c_sda_s1_readdata                          : std_logic_vector(31 downto 0); -- i2c_sda:readdata -> mm_interconnect_1:i2c_sda_s1_readdata
	signal mm_interconnect_1_i2c_sda_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_1:i2c_sda_s1_address -> i2c_sda:address
	signal mm_interconnect_1_i2c_sda_s1_write                             : std_logic;                     -- mm_interconnect_1:i2c_sda_s1_write -> mm_interconnect_1_i2c_sda_s1_write:in
	signal mm_interconnect_1_i2c_sda_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_1:i2c_sda_s1_writedata -> i2c_sda:writedata
	signal mm_interconnect_1_i2c_scl_s1_chipselect                        : std_logic;                     -- mm_interconnect_1:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	signal mm_interconnect_1_i2c_scl_s1_readdata                          : std_logic_vector(31 downto 0); -- i2c_scl:readdata -> mm_interconnect_1:i2c_scl_s1_readdata
	signal mm_interconnect_1_i2c_scl_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_1:i2c_scl_s1_address -> i2c_scl:address
	signal mm_interconnect_1_i2c_scl_s1_write                             : std_logic;                     -- mm_interconnect_1:i2c_scl_s1_write -> mm_interconnect_1_i2c_scl_s1_write:in
	signal mm_interconnect_1_i2c_scl_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_1:i2c_scl_s1_writedata -> i2c_scl:writedata
	signal mm_interconnect_1_ext_sensor_int_s1_chipselect                 : std_logic;                     -- mm_interconnect_1:ext_sensor_int_s1_chipselect -> ext_sensor_int:chipselect
	signal mm_interconnect_1_ext_sensor_int_s1_readdata                   : std_logic_vector(31 downto 0); -- ext_sensor_int:readdata -> mm_interconnect_1:ext_sensor_int_s1_readdata
	signal mm_interconnect_1_ext_sensor_int_s1_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_1:ext_sensor_int_s1_address -> ext_sensor_int:address
	signal mm_interconnect_1_ext_sensor_int_s1_write                      : std_logic;                     -- mm_interconnect_1:ext_sensor_int_s1_write -> mm_interconnect_1_ext_sensor_int_s1_write:in
	signal mm_interconnect_1_ext_sensor_int_s1_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_1:ext_sensor_int_s1_writedata -> ext_sensor_int:writedata
	signal mm_interconnect_1_i2c_ext_sda_s1_chipselect                    : std_logic;                     -- mm_interconnect_1:i2c_EXT_sda_s1_chipselect -> i2c_EXT_sda:chipselect
	signal mm_interconnect_1_i2c_ext_sda_s1_readdata                      : std_logic_vector(31 downto 0); -- i2c_EXT_sda:readdata -> mm_interconnect_1:i2c_EXT_sda_s1_readdata
	signal mm_interconnect_1_i2c_ext_sda_s1_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_1:i2c_EXT_sda_s1_address -> i2c_EXT_sda:address
	signal mm_interconnect_1_i2c_ext_sda_s1_write                         : std_logic;                     -- mm_interconnect_1:i2c_EXT_sda_s1_write -> mm_interconnect_1_i2c_ext_sda_s1_write:in
	signal mm_interconnect_1_i2c_ext_sda_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_1:i2c_EXT_sda_s1_writedata -> i2c_EXT_sda:writedata
	signal mm_interconnect_1_xbee_uart_s1_chipselect                      : std_logic;                     -- mm_interconnect_1:xbee_uart_s1_chipselect -> xbee_uart:chipselect
	signal mm_interconnect_1_xbee_uart_s1_readdata                        : std_logic_vector(15 downto 0); -- xbee_uart:readdata -> mm_interconnect_1:xbee_uart_s1_readdata
	signal mm_interconnect_1_xbee_uart_s1_address                         : std_logic_vector(2 downto 0);  -- mm_interconnect_1:xbee_uart_s1_address -> xbee_uart:address
	signal mm_interconnect_1_xbee_uart_s1_read                            : std_logic;                     -- mm_interconnect_1:xbee_uart_s1_read -> mm_interconnect_1_xbee_uart_s1_read:in
	signal mm_interconnect_1_xbee_uart_s1_begintransfer                   : std_logic;                     -- mm_interconnect_1:xbee_uart_s1_begintransfer -> xbee_uart:begintransfer
	signal mm_interconnect_1_xbee_uart_s1_write                           : std_logic;                     -- mm_interconnect_1:xbee_uart_s1_write -> mm_interconnect_1_xbee_uart_s1_write:in
	signal mm_interconnect_1_xbee_uart_s1_writedata                       : std_logic_vector(15 downto 0); -- mm_interconnect_1:xbee_uart_s1_writedata -> xbee_uart:writedata
	signal mm_interconnect_1_adc_spi_int_spi_control_port_chipselect      : std_logic;                     -- mm_interconnect_1:adc_spi_int_spi_control_port_chipselect -> adc_spi_int:spi_select
	signal mm_interconnect_1_adc_spi_int_spi_control_port_readdata        : std_logic_vector(15 downto 0); -- adc_spi_int:data_to_cpu -> mm_interconnect_1:adc_spi_int_spi_control_port_readdata
	signal mm_interconnect_1_adc_spi_int_spi_control_port_address         : std_logic_vector(2 downto 0);  -- mm_interconnect_1:adc_spi_int_spi_control_port_address -> adc_spi_int:mem_addr
	signal mm_interconnect_1_adc_spi_int_spi_control_port_read            : std_logic;                     -- mm_interconnect_1:adc_spi_int_spi_control_port_read -> mm_interconnect_1_adc_spi_int_spi_control_port_read:in
	signal mm_interconnect_1_adc_spi_int_spi_control_port_write           : std_logic;                     -- mm_interconnect_1:adc_spi_int_spi_control_port_write -> mm_interconnect_1_adc_spi_int_spi_control_port_write:in
	signal mm_interconnect_1_adc_spi_int_spi_control_port_writedata       : std_logic_vector(15 downto 0); -- mm_interconnect_1:adc_spi_int_spi_control_port_writedata -> adc_spi_int:data_from_cpu
	signal irq_mapper_receiver0_irq                                       : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal nios2_cpu_irq_irq                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_cpu:irq
	signal irq_mapper_receiver1_irq                                       : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	signal irq_synchronizer_receiver_irq                                  : std_logic_vector(0 downto 0);  -- epcs:irq -> irq_synchronizer:receiver_irq
	signal irq_mapper_receiver2_irq                                       : std_logic;                     -- irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	signal irq_synchronizer_001_receiver_irq                              : std_logic_vector(0 downto 0);  -- timer:irq -> irq_synchronizer_001:receiver_irq
	signal irq_mapper_receiver3_irq                                       : std_logic;                     -- irq_synchronizer_002:sender_irq -> irq_mapper:receiver3_irq
	signal irq_synchronizer_002_receiver_irq                              : std_logic_vector(0 downto 0);  -- pio_key:irq -> irq_synchronizer_002:receiver_irq
	signal irq_mapper_receiver4_irq                                       : std_logic;                     -- irq_synchronizer_003:sender_irq -> irq_mapper:receiver4_irq
	signal irq_synchronizer_003_receiver_irq                              : std_logic_vector(0 downto 0);  -- g_sensor_int:irq -> irq_synchronizer_003:receiver_irq
	signal irq_mapper_receiver5_irq                                       : std_logic;                     -- irq_synchronizer_004:sender_irq -> irq_mapper:receiver5_irq
	signal irq_synchronizer_004_receiver_irq                              : std_logic_vector(0 downto 0);  -- ext_sensor_int:irq -> irq_synchronizer_004:receiver_irq
	signal irq_mapper_receiver6_irq                                       : std_logic;                     -- irq_synchronizer_005:sender_irq -> irq_mapper:receiver6_irq
	signal irq_synchronizer_005_receiver_irq                              : std_logic_vector(0 downto 0);  -- adc_spi_int:irq -> irq_synchronizer_005:receiver_irq
	signal irq_mapper_receiver7_irq                                       : std_logic;                     -- irq_synchronizer_006:sender_irq -> irq_mapper:receiver7_irq
	signal irq_synchronizer_006_receiver_irq                              : std_logic_vector(0 downto 0);  -- xbee_uart:irq -> irq_synchronizer_006:receiver_irq
	signal rst_controller_reset_out_reset                                 : std_logic;                     -- rst_controller:reset_out -> [clock_crossing_bridge_IO:m0_reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, irq_synchronizer_005:receiver_reset, irq_synchronizer_006:receiver_reset, mm_interconnect_1:clock_crossing_bridge_IO_m0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                             : std_logic;                     -- rst_controller:reset_req -> [epcs:reset_req, rst_translator:reset_req_in]
	signal nios2_cpu_debug_reset_request_reset                            : std_logic;                     -- nios2_cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in0, rst_controller_002:reset_in1]
	signal rst_controller_001_reset_out_reset                             : std_logic;                     -- rst_controller_001:reset_out -> [altpll_sys:reset, mm_interconnect_0:altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal rst_controller_002_reset_out_reset                             : std_logic;                     -- rst_controller_002:reset_out -> [clock_crossing_bridge_IO:s0_reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, irq_synchronizer_005:sender_reset, irq_synchronizer_006:sender_reset, mm_interconnect_0:nios2_cpu_reset_reset_bridge_in_reset_reset, onchip_mem:reset, rst_controller_002_reset_out_reset:in, rst_translator_001:in_reset]
	signal rst_controller_002_reset_out_reset_req                         : std_logic;                     -- rst_controller_002:reset_req -> [nios2_cpu:reset_req, onchip_mem:reset_req, rst_translator_001:reset_req_in]
	signal reset_reset_n_ports_inv                                        : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv   : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                      : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_1_epcs_epcs_control_port_read_ports_inv        : std_logic;                     -- mm_interconnect_1_epcs_epcs_control_port_read:inv -> epcs:read_n
	signal mm_interconnect_1_epcs_epcs_control_port_write_ports_inv       : std_logic;                     -- mm_interconnect_1_epcs_epcs_control_port_write:inv -> epcs:write_n
	signal mm_interconnect_1_timer_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_1_timer_s1_write:inv -> timer:write_n
	signal mm_interconnect_1_pio_leds_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_1_pio_leds_s1_write:inv -> pio_leds:write_n
	signal mm_interconnect_1_pio_key_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_1_pio_key_s1_write:inv -> pio_key:write_n
	signal mm_interconnect_1_g_sensor_int_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_1_g_sensor_int_s1_write:inv -> g_sensor_int:write_n
	signal mm_interconnect_1_i2c_sda_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_1_i2c_sda_s1_write:inv -> i2c_sda:write_n
	signal mm_interconnect_1_i2c_scl_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_1_i2c_scl_s1_write:inv -> i2c_scl:write_n
	signal mm_interconnect_1_ext_sensor_int_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_1_ext_sensor_int_s1_write:inv -> ext_sensor_int:write_n
	signal mm_interconnect_1_i2c_ext_sda_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_1_i2c_ext_sda_s1_write:inv -> i2c_EXT_sda:write_n
	signal mm_interconnect_1_xbee_uart_s1_read_ports_inv                  : std_logic;                     -- mm_interconnect_1_xbee_uart_s1_read:inv -> xbee_uart:read_n
	signal mm_interconnect_1_xbee_uart_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_1_xbee_uart_s1_write:inv -> xbee_uart:write_n
	signal mm_interconnect_1_adc_spi_int_spi_control_port_read_ports_inv  : std_logic;                     -- mm_interconnect_1_adc_spi_int_spi_control_port_read:inv -> adc_spi_int:read_n
	signal mm_interconnect_1_adc_spi_int_spi_control_port_write_ports_inv : std_logic;                     -- mm_interconnect_1_adc_spi_int_spi_control_port_write:inv -> adc_spi_int:write_n
	signal rst_controller_reset_out_reset_ports_inv                       : std_logic;                     -- rst_controller_reset_out_reset:inv -> [adc_spi_int:reset_n, epcs:reset_n, ext_sensor_int:reset_n, g_sensor_int:reset_n, i2c_EXT_sda:reset_n, i2c_scl:reset_n, i2c_sda:reset_n, pio_key:reset_n, pio_leds:reset_n, pio_switch:reset_n, sysid_qsys:reset_n, timer:reset_n, xbee_uart:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                   : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> [jtag_uart:rst_n, nios2_cpu:reset_n, sdram:reset_n]

begin

	adc_spi_int : component DE0_nano_system_adc_spi_int
		port map (
			clk           => altpll_sys_c2_clk,                                              --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                       --            reset.reset_n
			data_from_cpu => mm_interconnect_1_adc_spi_int_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_1_adc_spi_int_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_1_adc_spi_int_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_1_adc_spi_int_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_1_adc_spi_int_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_1_adc_spi_int_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_synchronizer_005_receiver_irq(0),                           --              irq.irq
			MISO          => adc_spi_conduit_MISO,                                           --         external.export
			MOSI          => adc_spi_conduit_MOSI,                                           --                 .export
			SCLK          => adc_spi_conduit_SCLK,                                           --                 .export
			SS_n          => adc_spi_conduit_SS_n                                            --                 .export
		);

	altpll_sys : component DE0_nano_system_altpll_sys
		port map (
			clk                => clk_clk,                                          --       inclk_interface.clk
			reset              => rst_controller_001_reset_out_reset,               -- inclk_interface_reset.reset
			read               => mm_interconnect_0_altpll_sys_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_altpll_sys_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_altpll_sys_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_altpll_sys_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_altpll_sys_pll_slave_writedata, --                      .writedata
			c0                 => altpll_sys_c0_clk,                                --                    c0.clk
			c1                 => altpll_sys_c1_clk,                                --                    c1.clk
			c2                 => altpll_sys_c2_clk,                                --                    c2.clk
			locked             => altpll_sys_locked_conduit_export,                 --        locked_conduit.export
			scandone           => open,                                             --           (terminated)
			scandataout        => open,                                             --           (terminated)
			phasecounterselect => "0000",                                           --           (terminated)
			phaseupdown        => '0',                                              --           (terminated)
			phasestep          => '0',                                              --           (terminated)
			scanclk            => '0',                                              --           (terminated)
			scanclkena         => '0',                                              --           (terminated)
			scandata           => '0',                                              --           (terminated)
			configupdate       => '0',                                              --           (terminated)
			areset             => '0',                                              --           (terminated)
			phasedone          => open                                              --           (terminated)
		);

	clock_crossing_bridge_io : component altera_avalon_mm_clock_crossing_bridge
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			HDL_ADDR_WIDTH      => 12,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 16,
			RESPONSE_FIFO_DEPTH => 32,
			MASTER_SYNC_DEPTH   => 3,
			SLAVE_SYNC_DEPTH    => 3
		)
		port map (
			m0_clk           => altpll_sys_c2_clk,                                           --   m0_clk.clk
			m0_reset         => rst_controller_reset_out_reset,                              -- m0_reset.reset
			s0_clk           => altpll_sys_c0_clk,                                           --   s0_clk.clk
			s0_reset         => rst_controller_002_reset_out_reset,                          -- s0_reset.reset
			s0_waitrequest   => mm_interconnect_0_clock_crossing_bridge_io_s0_waitrequest,   --       s0.waitrequest
			s0_readdata      => mm_interconnect_0_clock_crossing_bridge_io_s0_readdata,      --         .readdata
			s0_readdatavalid => mm_interconnect_0_clock_crossing_bridge_io_s0_readdatavalid, --         .readdatavalid
			s0_burstcount    => mm_interconnect_0_clock_crossing_bridge_io_s0_burstcount,    --         .burstcount
			s0_writedata     => mm_interconnect_0_clock_crossing_bridge_io_s0_writedata,     --         .writedata
			s0_address       => mm_interconnect_0_clock_crossing_bridge_io_s0_address,       --         .address
			s0_write         => mm_interconnect_0_clock_crossing_bridge_io_s0_write,         --         .write
			s0_read          => mm_interconnect_0_clock_crossing_bridge_io_s0_read,          --         .read
			s0_byteenable    => mm_interconnect_0_clock_crossing_bridge_io_s0_byteenable,    --         .byteenable
			s0_debugaccess   => mm_interconnect_0_clock_crossing_bridge_io_s0_debugaccess,   --         .debugaccess
			m0_waitrequest   => clock_crossing_bridge_io_m0_waitrequest,                     --       m0.waitrequest
			m0_readdata      => clock_crossing_bridge_io_m0_readdata,                        --         .readdata
			m0_readdatavalid => clock_crossing_bridge_io_m0_readdatavalid,                   --         .readdatavalid
			m0_burstcount    => clock_crossing_bridge_io_m0_burstcount,                      --         .burstcount
			m0_writedata     => clock_crossing_bridge_io_m0_writedata,                       --         .writedata
			m0_address       => clock_crossing_bridge_io_m0_address,                         --         .address
			m0_write         => clock_crossing_bridge_io_m0_write,                           --         .write
			m0_read          => clock_crossing_bridge_io_m0_read,                            --         .read
			m0_byteenable    => clock_crossing_bridge_io_m0_byteenable,                      --         .byteenable
			m0_debugaccess   => clock_crossing_bridge_io_m0_debugaccess                      --         .debugaccess
		);

	epcs : component DE0_nano_system_epcs
		port map (
			clk        => altpll_sys_c2_clk,                                        --               clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                 --             reset.reset_n
			reset_req  => rst_controller_reset_out_reset_req,                       --                  .reset_req
			address    => mm_interconnect_1_epcs_epcs_control_port_address,         -- epcs_control_port.address
			chipselect => mm_interconnect_1_epcs_epcs_control_port_chipselect,      --                  .chipselect
			read_n     => mm_interconnect_1_epcs_epcs_control_port_read_ports_inv,  --                  .read_n
			readdata   => mm_interconnect_1_epcs_epcs_control_port_readdata,        --                  .readdata
			write_n    => mm_interconnect_1_epcs_epcs_control_port_write_ports_inv, --                  .write_n
			writedata  => mm_interconnect_1_epcs_epcs_control_port_writedata,       --                  .writedata
			irq        => irq_synchronizer_receiver_irq(0),                         --               irq.irq
			dclk       => epcs_dclk,                                                --          external.export
			sce        => epcs_sce,                                                 --                  .export
			sdo        => epcs_sdo,                                                 --                  .export
			data0      => epcs_data0                                                --                  .export
		);

	ext_sensor_int : component DE0_nano_system_ext_sensor_int
		port map (
			clk        => altpll_sys_c2_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address    => mm_interconnect_1_ext_sensor_int_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_ext_sensor_int_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_ext_sensor_int_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_ext_sensor_int_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_ext_sensor_int_s1_readdata,        --                    .readdata
			in_port    => ext_sensor_irq_export,                               -- external_connection.export
			irq        => irq_synchronizer_004_receiver_irq(0)                 --                 irq.irq
		);

	g_sensor_int : component DE0_nano_system_g_sensor_int
		port map (
			clk        => altpll_sys_c2_clk,                                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_1_g_sensor_int_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_g_sensor_int_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_g_sensor_int_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_g_sensor_int_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_g_sensor_int_s1_readdata,        --                    .readdata
			in_port    => g_sensor_irq_export,                               -- external_connection.export
			irq        => irq_synchronizer_003_receiver_irq(0)               --                 irq.irq
		);

	i2c_ext_sda : component DE0_nano_system_i2c_EXT_sda
		port map (
			clk        => altpll_sys_c2_clk,                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_1_i2c_ext_sda_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_i2c_ext_sda_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_i2c_ext_sda_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_i2c_ext_sda_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_i2c_ext_sda_s1_readdata,        --                    .readdata
			bidir_port => i2c_ext_sda_export                                -- external_connection.export
		);

	i2c_scl : component DE0_nano_system_i2c_scl
		port map (
			clk        => altpll_sys_c2_clk,                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_1_i2c_scl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_i2c_scl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_i2c_scl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_i2c_scl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_i2c_scl_s1_readdata,        --                    .readdata
			out_port   => i2c_scl_export                                -- external_connection.export
		);

	i2c_sda : component DE0_nano_system_i2c_EXT_sda
		port map (
			clk        => altpll_sys_c2_clk,                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_1_i2c_sda_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_i2c_sda_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_i2c_sda_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_i2c_sda_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_i2c_sda_s1_readdata,        --                    .readdata
			bidir_port => i2c_sda_export                                -- external_connection.export
		);

	jtag_uart : component DE0_nano_system_jtag_uart
		port map (
			clk            => altpll_sys_c0_clk,                                             --               clk.clk
			rst_n          => rst_controller_002_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	nios2_cpu : component DE0_nano_system_nios2_cpu
		port map (
			clk                                 => altpll_sys_c0_clk,                                       --                       clk.clk
			reset_n                             => rst_controller_002_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_002_reset_out_reset_req,                  --                          .reset_req
			d_address                           => nios2_cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_cpu_data_master_read,                              --                          .read
			d_readdata                          => nios2_cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_cpu_data_master_write,                             --                          .write
			d_writedata                         => nios2_cpu_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_cpu_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_cpu_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                     -- custom_instruction_master.readra
		);

	onchip_mem : component DE0_nano_system_onchip_mem
		port map (
			clk        => altpll_sys_c0_clk,                          --   clk1.clk
			address    => mm_interconnect_0_onchip_mem_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_mem_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_mem_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_mem_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_mem_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_mem_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_mem_s1_byteenable, --       .byteenable
			reset      => rst_controller_002_reset_out_reset,         -- reset1.reset
			reset_req  => rst_controller_002_reset_out_reset_req,     --       .reset_req
			freeze     => '0'                                         -- (terminated)
		);

	pio_key : component DE0_nano_system_pio_key
		port map (
			clk        => altpll_sys_c2_clk,                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_1_pio_key_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_pio_key_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_pio_key_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_pio_key_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_pio_key_s1_readdata,        --                    .readdata
			in_port    => pio_key_export,                               -- external_connection.export
			irq        => irq_synchronizer_002_receiver_irq(0)          --                 irq.irq
		);

	pio_leds : component DE0_nano_system_pio_leds
		port map (
			clk        => altpll_sys_c2_clk,                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_1_pio_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_pio_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_pio_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_pio_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_pio_leds_s1_readdata,        --                    .readdata
			out_port   => pio_leds_export                                -- external_connection.export
		);

	pio_switch : component DE0_nano_system_pio_switch
		port map (
			clk      => altpll_sys_c2_clk,                        --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_1_pio_switch_s1_address,  --                  s1.address
			readdata => mm_interconnect_1_pio_switch_s1_readdata, --                    .readdata
			in_port  => pio_switch_export                         -- external_connection.export
		);

	sdram : component DE0_nano_system_sdram
		port map (
			clk            => altpll_sys_c0_clk,                               --   clk.clk
			reset_n        => rst_controller_002_reset_out_reset_ports_inv,    -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	sysid_qsys : component DE0_nano_system_sysid_qsys
		port map (
			clock    => altpll_sys_c2_clk,                                     --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,              --         reset.reset_n
			readdata => mm_interconnect_1_sysid_qsys_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_1_sysid_qsys_control_slave_address(0)  --              .address
		);

	timer : component DE0_nano_system_timer
		port map (
			clk        => altpll_sys_c2_clk,                          --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   -- reset.reset_n
			address    => mm_interconnect_1_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_1_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_1_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_1_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_1_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_synchronizer_001_receiver_irq(0)        --   irq.irq
		);

	xbee_uart : component DE0_nano_system_xbee_uart
		port map (
			clk           => altpll_sys_c2_clk,                              --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address       => mm_interconnect_1_xbee_uart_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_1_xbee_uart_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_1_xbee_uart_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_1_xbee_uart_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_1_xbee_uart_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_1_xbee_uart_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_1_xbee_uart_s1_readdata,        --                    .readdata
			rxd           => xbee_rxd,                                       -- external_connection.export
			txd           => xbee_txd,                                       --                    .export
			irq           => irq_synchronizer_006_receiver_irq(0)            --                 irq.irq
		);

	mm_interconnect_0 : component DE0_nano_system_mm_interconnect_0
		port map (
			altpll_sys_c0_clk                                            => altpll_sys_c0_clk,                                           --                                          altpll_sys_c0.clk
			clk_50_clk_clk                                               => clk_clk,                                                     --                                             clk_50_clk.clk
			altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                          -- altpll_sys_inclk_interface_reset_reset_bridge_in_reset.reset
			nios2_cpu_reset_reset_bridge_in_reset_reset                  => rst_controller_002_reset_out_reset,                          --                  nios2_cpu_reset_reset_bridge_in_reset.reset
			nios2_cpu_data_master_address                                => nios2_cpu_data_master_address,                               --                                  nios2_cpu_data_master.address
			nios2_cpu_data_master_waitrequest                            => nios2_cpu_data_master_waitrequest,                           --                                                       .waitrequest
			nios2_cpu_data_master_byteenable                             => nios2_cpu_data_master_byteenable,                            --                                                       .byteenable
			nios2_cpu_data_master_read                                   => nios2_cpu_data_master_read,                                  --                                                       .read
			nios2_cpu_data_master_readdata                               => nios2_cpu_data_master_readdata,                              --                                                       .readdata
			nios2_cpu_data_master_readdatavalid                          => nios2_cpu_data_master_readdatavalid,                         --                                                       .readdatavalid
			nios2_cpu_data_master_write                                  => nios2_cpu_data_master_write,                                 --                                                       .write
			nios2_cpu_data_master_writedata                              => nios2_cpu_data_master_writedata,                             --                                                       .writedata
			nios2_cpu_data_master_debugaccess                            => nios2_cpu_data_master_debugaccess,                           --                                                       .debugaccess
			nios2_cpu_instruction_master_address                         => nios2_cpu_instruction_master_address,                        --                           nios2_cpu_instruction_master.address
			nios2_cpu_instruction_master_waitrequest                     => nios2_cpu_instruction_master_waitrequest,                    --                                                       .waitrequest
			nios2_cpu_instruction_master_read                            => nios2_cpu_instruction_master_read,                           --                                                       .read
			nios2_cpu_instruction_master_readdata                        => nios2_cpu_instruction_master_readdata,                       --                                                       .readdata
			nios2_cpu_instruction_master_readdatavalid                   => nios2_cpu_instruction_master_readdatavalid,                  --                                                       .readdatavalid
			altpll_sys_pll_slave_address                                 => mm_interconnect_0_altpll_sys_pll_slave_address,              --                                   altpll_sys_pll_slave.address
			altpll_sys_pll_slave_write                                   => mm_interconnect_0_altpll_sys_pll_slave_write,                --                                                       .write
			altpll_sys_pll_slave_read                                    => mm_interconnect_0_altpll_sys_pll_slave_read,                 --                                                       .read
			altpll_sys_pll_slave_readdata                                => mm_interconnect_0_altpll_sys_pll_slave_readdata,             --                                                       .readdata
			altpll_sys_pll_slave_writedata                               => mm_interconnect_0_altpll_sys_pll_slave_writedata,            --                                                       .writedata
			clock_crossing_bridge_IO_s0_address                          => mm_interconnect_0_clock_crossing_bridge_io_s0_address,       --                            clock_crossing_bridge_IO_s0.address
			clock_crossing_bridge_IO_s0_write                            => mm_interconnect_0_clock_crossing_bridge_io_s0_write,         --                                                       .write
			clock_crossing_bridge_IO_s0_read                             => mm_interconnect_0_clock_crossing_bridge_io_s0_read,          --                                                       .read
			clock_crossing_bridge_IO_s0_readdata                         => mm_interconnect_0_clock_crossing_bridge_io_s0_readdata,      --                                                       .readdata
			clock_crossing_bridge_IO_s0_writedata                        => mm_interconnect_0_clock_crossing_bridge_io_s0_writedata,     --                                                       .writedata
			clock_crossing_bridge_IO_s0_burstcount                       => mm_interconnect_0_clock_crossing_bridge_io_s0_burstcount,    --                                                       .burstcount
			clock_crossing_bridge_IO_s0_byteenable                       => mm_interconnect_0_clock_crossing_bridge_io_s0_byteenable,    --                                                       .byteenable
			clock_crossing_bridge_IO_s0_readdatavalid                    => mm_interconnect_0_clock_crossing_bridge_io_s0_readdatavalid, --                                                       .readdatavalid
			clock_crossing_bridge_IO_s0_waitrequest                      => mm_interconnect_0_clock_crossing_bridge_io_s0_waitrequest,   --                                                       .waitrequest
			clock_crossing_bridge_IO_s0_debugaccess                      => mm_interconnect_0_clock_crossing_bridge_io_s0_debugaccess,   --                                                       .debugaccess
			jtag_uart_avalon_jtag_slave_address                          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,       --                            jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                            => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,         --                                                       .write
			jtag_uart_avalon_jtag_slave_read                             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,          --                                                       .read
			jtag_uart_avalon_jtag_slave_readdata                         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,      --                                                       .readdata
			jtag_uart_avalon_jtag_slave_writedata                        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,     --                                                       .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,   --                                                       .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,    --                                                       .chipselect
			nios2_cpu_debug_mem_slave_address                            => mm_interconnect_0_nios2_cpu_debug_mem_slave_address,         --                              nios2_cpu_debug_mem_slave.address
			nios2_cpu_debug_mem_slave_write                              => mm_interconnect_0_nios2_cpu_debug_mem_slave_write,           --                                                       .write
			nios2_cpu_debug_mem_slave_read                               => mm_interconnect_0_nios2_cpu_debug_mem_slave_read,            --                                                       .read
			nios2_cpu_debug_mem_slave_readdata                           => mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata,        --                                                       .readdata
			nios2_cpu_debug_mem_slave_writedata                          => mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata,       --                                                       .writedata
			nios2_cpu_debug_mem_slave_byteenable                         => mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable,      --                                                       .byteenable
			nios2_cpu_debug_mem_slave_waitrequest                        => mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest,     --                                                       .waitrequest
			nios2_cpu_debug_mem_slave_debugaccess                        => mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess,     --                                                       .debugaccess
			onchip_mem_s1_address                                        => mm_interconnect_0_onchip_mem_s1_address,                     --                                          onchip_mem_s1.address
			onchip_mem_s1_write                                          => mm_interconnect_0_onchip_mem_s1_write,                       --                                                       .write
			onchip_mem_s1_readdata                                       => mm_interconnect_0_onchip_mem_s1_readdata,                    --                                                       .readdata
			onchip_mem_s1_writedata                                      => mm_interconnect_0_onchip_mem_s1_writedata,                   --                                                       .writedata
			onchip_mem_s1_byteenable                                     => mm_interconnect_0_onchip_mem_s1_byteenable,                  --                                                       .byteenable
			onchip_mem_s1_chipselect                                     => mm_interconnect_0_onchip_mem_s1_chipselect,                  --                                                       .chipselect
			onchip_mem_s1_clken                                          => mm_interconnect_0_onchip_mem_s1_clken,                       --                                                       .clken
			sdram_s1_address                                             => mm_interconnect_0_sdram_s1_address,                          --                                               sdram_s1.address
			sdram_s1_write                                               => mm_interconnect_0_sdram_s1_write,                            --                                                       .write
			sdram_s1_read                                                => mm_interconnect_0_sdram_s1_read,                             --                                                       .read
			sdram_s1_readdata                                            => mm_interconnect_0_sdram_s1_readdata,                         --                                                       .readdata
			sdram_s1_writedata                                           => mm_interconnect_0_sdram_s1_writedata,                        --                                                       .writedata
			sdram_s1_byteenable                                          => mm_interconnect_0_sdram_s1_byteenable,                       --                                                       .byteenable
			sdram_s1_readdatavalid                                       => mm_interconnect_0_sdram_s1_readdatavalid,                    --                                                       .readdatavalid
			sdram_s1_waitrequest                                         => mm_interconnect_0_sdram_s1_waitrequest,                      --                                                       .waitrequest
			sdram_s1_chipselect                                          => mm_interconnect_0_sdram_s1_chipselect                        --                                                       .chipselect
		);

	mm_interconnect_1 : component DE0_nano_system_mm_interconnect_1
		port map (
			altpll_sys_c2_clk                                             => altpll_sys_c2_clk,                                         --                                           altpll_sys_c2.clk
			clock_crossing_bridge_IO_m0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- clock_crossing_bridge_IO_m0_reset_reset_bridge_in_reset.reset
			clock_crossing_bridge_IO_m0_address                           => clock_crossing_bridge_io_m0_address,                       --                             clock_crossing_bridge_IO_m0.address
			clock_crossing_bridge_IO_m0_waitrequest                       => clock_crossing_bridge_io_m0_waitrequest,                   --                                                        .waitrequest
			clock_crossing_bridge_IO_m0_burstcount                        => clock_crossing_bridge_io_m0_burstcount,                    --                                                        .burstcount
			clock_crossing_bridge_IO_m0_byteenable                        => clock_crossing_bridge_io_m0_byteenable,                    --                                                        .byteenable
			clock_crossing_bridge_IO_m0_read                              => clock_crossing_bridge_io_m0_read,                          --                                                        .read
			clock_crossing_bridge_IO_m0_readdata                          => clock_crossing_bridge_io_m0_readdata,                      --                                                        .readdata
			clock_crossing_bridge_IO_m0_readdatavalid                     => clock_crossing_bridge_io_m0_readdatavalid,                 --                                                        .readdatavalid
			clock_crossing_bridge_IO_m0_write                             => clock_crossing_bridge_io_m0_write,                         --                                                        .write
			clock_crossing_bridge_IO_m0_writedata                         => clock_crossing_bridge_io_m0_writedata,                     --                                                        .writedata
			clock_crossing_bridge_IO_m0_debugaccess                       => clock_crossing_bridge_io_m0_debugaccess,                   --                                                        .debugaccess
			adc_spi_int_spi_control_port_address                          => mm_interconnect_1_adc_spi_int_spi_control_port_address,    --                            adc_spi_int_spi_control_port.address
			adc_spi_int_spi_control_port_write                            => mm_interconnect_1_adc_spi_int_spi_control_port_write,      --                                                        .write
			adc_spi_int_spi_control_port_read                             => mm_interconnect_1_adc_spi_int_spi_control_port_read,       --                                                        .read
			adc_spi_int_spi_control_port_readdata                         => mm_interconnect_1_adc_spi_int_spi_control_port_readdata,   --                                                        .readdata
			adc_spi_int_spi_control_port_writedata                        => mm_interconnect_1_adc_spi_int_spi_control_port_writedata,  --                                                        .writedata
			adc_spi_int_spi_control_port_chipselect                       => mm_interconnect_1_adc_spi_int_spi_control_port_chipselect, --                                                        .chipselect
			epcs_epcs_control_port_address                                => mm_interconnect_1_epcs_epcs_control_port_address,          --                                  epcs_epcs_control_port.address
			epcs_epcs_control_port_write                                  => mm_interconnect_1_epcs_epcs_control_port_write,            --                                                        .write
			epcs_epcs_control_port_read                                   => mm_interconnect_1_epcs_epcs_control_port_read,             --                                                        .read
			epcs_epcs_control_port_readdata                               => mm_interconnect_1_epcs_epcs_control_port_readdata,         --                                                        .readdata
			epcs_epcs_control_port_writedata                              => mm_interconnect_1_epcs_epcs_control_port_writedata,        --                                                        .writedata
			epcs_epcs_control_port_chipselect                             => mm_interconnect_1_epcs_epcs_control_port_chipselect,       --                                                        .chipselect
			ext_sensor_int_s1_address                                     => mm_interconnect_1_ext_sensor_int_s1_address,               --                                       ext_sensor_int_s1.address
			ext_sensor_int_s1_write                                       => mm_interconnect_1_ext_sensor_int_s1_write,                 --                                                        .write
			ext_sensor_int_s1_readdata                                    => mm_interconnect_1_ext_sensor_int_s1_readdata,              --                                                        .readdata
			ext_sensor_int_s1_writedata                                   => mm_interconnect_1_ext_sensor_int_s1_writedata,             --                                                        .writedata
			ext_sensor_int_s1_chipselect                                  => mm_interconnect_1_ext_sensor_int_s1_chipselect,            --                                                        .chipselect
			g_sensor_int_s1_address                                       => mm_interconnect_1_g_sensor_int_s1_address,                 --                                         g_sensor_int_s1.address
			g_sensor_int_s1_write                                         => mm_interconnect_1_g_sensor_int_s1_write,                   --                                                        .write
			g_sensor_int_s1_readdata                                      => mm_interconnect_1_g_sensor_int_s1_readdata,                --                                                        .readdata
			g_sensor_int_s1_writedata                                     => mm_interconnect_1_g_sensor_int_s1_writedata,               --                                                        .writedata
			g_sensor_int_s1_chipselect                                    => mm_interconnect_1_g_sensor_int_s1_chipselect,              --                                                        .chipselect
			i2c_EXT_sda_s1_address                                        => mm_interconnect_1_i2c_ext_sda_s1_address,                  --                                          i2c_EXT_sda_s1.address
			i2c_EXT_sda_s1_write                                          => mm_interconnect_1_i2c_ext_sda_s1_write,                    --                                                        .write
			i2c_EXT_sda_s1_readdata                                       => mm_interconnect_1_i2c_ext_sda_s1_readdata,                 --                                                        .readdata
			i2c_EXT_sda_s1_writedata                                      => mm_interconnect_1_i2c_ext_sda_s1_writedata,                --                                                        .writedata
			i2c_EXT_sda_s1_chipselect                                     => mm_interconnect_1_i2c_ext_sda_s1_chipselect,               --                                                        .chipselect
			i2c_scl_s1_address                                            => mm_interconnect_1_i2c_scl_s1_address,                      --                                              i2c_scl_s1.address
			i2c_scl_s1_write                                              => mm_interconnect_1_i2c_scl_s1_write,                        --                                                        .write
			i2c_scl_s1_readdata                                           => mm_interconnect_1_i2c_scl_s1_readdata,                     --                                                        .readdata
			i2c_scl_s1_writedata                                          => mm_interconnect_1_i2c_scl_s1_writedata,                    --                                                        .writedata
			i2c_scl_s1_chipselect                                         => mm_interconnect_1_i2c_scl_s1_chipselect,                   --                                                        .chipselect
			i2c_sda_s1_address                                            => mm_interconnect_1_i2c_sda_s1_address,                      --                                              i2c_sda_s1.address
			i2c_sda_s1_write                                              => mm_interconnect_1_i2c_sda_s1_write,                        --                                                        .write
			i2c_sda_s1_readdata                                           => mm_interconnect_1_i2c_sda_s1_readdata,                     --                                                        .readdata
			i2c_sda_s1_writedata                                          => mm_interconnect_1_i2c_sda_s1_writedata,                    --                                                        .writedata
			i2c_sda_s1_chipselect                                         => mm_interconnect_1_i2c_sda_s1_chipselect,                   --                                                        .chipselect
			pio_key_s1_address                                            => mm_interconnect_1_pio_key_s1_address,                      --                                              pio_key_s1.address
			pio_key_s1_write                                              => mm_interconnect_1_pio_key_s1_write,                        --                                                        .write
			pio_key_s1_readdata                                           => mm_interconnect_1_pio_key_s1_readdata,                     --                                                        .readdata
			pio_key_s1_writedata                                          => mm_interconnect_1_pio_key_s1_writedata,                    --                                                        .writedata
			pio_key_s1_chipselect                                         => mm_interconnect_1_pio_key_s1_chipselect,                   --                                                        .chipselect
			pio_leds_s1_address                                           => mm_interconnect_1_pio_leds_s1_address,                     --                                             pio_leds_s1.address
			pio_leds_s1_write                                             => mm_interconnect_1_pio_leds_s1_write,                       --                                                        .write
			pio_leds_s1_readdata                                          => mm_interconnect_1_pio_leds_s1_readdata,                    --                                                        .readdata
			pio_leds_s1_writedata                                         => mm_interconnect_1_pio_leds_s1_writedata,                   --                                                        .writedata
			pio_leds_s1_chipselect                                        => mm_interconnect_1_pio_leds_s1_chipselect,                  --                                                        .chipselect
			pio_switch_s1_address                                         => mm_interconnect_1_pio_switch_s1_address,                   --                                           pio_switch_s1.address
			pio_switch_s1_readdata                                        => mm_interconnect_1_pio_switch_s1_readdata,                  --                                                        .readdata
			sysid_qsys_control_slave_address                              => mm_interconnect_1_sysid_qsys_control_slave_address,        --                                sysid_qsys_control_slave.address
			sysid_qsys_control_slave_readdata                             => mm_interconnect_1_sysid_qsys_control_slave_readdata,       --                                                        .readdata
			timer_s1_address                                              => mm_interconnect_1_timer_s1_address,                        --                                                timer_s1.address
			timer_s1_write                                                => mm_interconnect_1_timer_s1_write,                          --                                                        .write
			timer_s1_readdata                                             => mm_interconnect_1_timer_s1_readdata,                       --                                                        .readdata
			timer_s1_writedata                                            => mm_interconnect_1_timer_s1_writedata,                      --                                                        .writedata
			timer_s1_chipselect                                           => mm_interconnect_1_timer_s1_chipselect,                     --                                                        .chipselect
			xbee_uart_s1_address                                          => mm_interconnect_1_xbee_uart_s1_address,                    --                                            xbee_uart_s1.address
			xbee_uart_s1_write                                            => mm_interconnect_1_xbee_uart_s1_write,                      --                                                        .write
			xbee_uart_s1_read                                             => mm_interconnect_1_xbee_uart_s1_read,                       --                                                        .read
			xbee_uart_s1_readdata                                         => mm_interconnect_1_xbee_uart_s1_readdata,                   --                                                        .readdata
			xbee_uart_s1_writedata                                        => mm_interconnect_1_xbee_uart_s1_writedata,                  --                                                        .writedata
			xbee_uart_s1_begintransfer                                    => mm_interconnect_1_xbee_uart_s1_begintransfer,              --                                                        .begintransfer
			xbee_uart_s1_chipselect                                       => mm_interconnect_1_xbee_uart_s1_chipselect                  --                                                        .chipselect
		);

	irq_mapper : component DE0_nano_system_irq_mapper
		port map (
			clk           => altpll_sys_c0_clk,                  --       clk.clk
			reset         => rst_controller_002_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,           -- receiver5.irq
			receiver6_irq => irq_mapper_receiver6_irq,           -- receiver6.irq
			receiver7_irq => irq_mapper_receiver7_irq,           -- receiver7.irq
			sender_irq    => nios2_cpu_irq_irq                   --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => altpll_sys_c2_clk,                  --       receiver_clk.clk
			sender_clk     => altpll_sys_c0_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_002_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver1_irq            --             sender.irq
		);

	irq_synchronizer_001 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => altpll_sys_c2_clk,                  --       receiver_clk.clk
			sender_clk     => altpll_sys_c0_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_002_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_001_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver2_irq            --             sender.irq
		);

	irq_synchronizer_002 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => altpll_sys_c2_clk,                  --       receiver_clk.clk
			sender_clk     => altpll_sys_c0_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_002_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_002_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver3_irq            --             sender.irq
		);

	irq_synchronizer_003 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => altpll_sys_c2_clk,                  --       receiver_clk.clk
			sender_clk     => altpll_sys_c0_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_002_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_003_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver4_irq            --             sender.irq
		);

	irq_synchronizer_004 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => altpll_sys_c2_clk,                  --       receiver_clk.clk
			sender_clk     => altpll_sys_c0_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_002_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_004_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver5_irq            --             sender.irq
		);

	irq_synchronizer_005 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => altpll_sys_c2_clk,                  --       receiver_clk.clk
			sender_clk     => altpll_sys_c0_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_002_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_005_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver6_irq            --             sender.irq
		);

	irq_synchronizer_006 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => altpll_sys_c2_clk,                  --       receiver_clk.clk
			sender_clk     => altpll_sys_c0_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_002_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_006_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver7_irq            --             sender.irq
		);

	rst_controller : component de0_nano_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,             -- reset_in0.reset
			reset_in1      => nios2_cpu_debug_reset_request_reset, -- reset_in1.reset
			clk            => altpll_sys_c2_clk,                   --       clk.clk
			reset_out      => rst_controller_reset_out_reset,      -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,  --          .reset_req
			reset_req_in0  => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_in2      => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	rst_controller_001 : component de0_nano_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_cpu_debug_reset_request_reset, -- reset_in0.reset
			clk            => clk_clk,                             --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,  -- reset_out.reset
			reset_req      => open,                                -- (terminated)
			reset_req_in0  => '0',                                 -- (terminated)
			reset_in1      => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_in2      => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	rst_controller_002 : component de0_nano_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_cpu_debug_reset_request_reset,    -- reset_in1.reset
			clk            => altpll_sys_c0_clk,                      --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_1_epcs_epcs_control_port_read_ports_inv <= not mm_interconnect_1_epcs_epcs_control_port_read;

	mm_interconnect_1_epcs_epcs_control_port_write_ports_inv <= not mm_interconnect_1_epcs_epcs_control_port_write;

	mm_interconnect_1_timer_s1_write_ports_inv <= not mm_interconnect_1_timer_s1_write;

	mm_interconnect_1_pio_leds_s1_write_ports_inv <= not mm_interconnect_1_pio_leds_s1_write;

	mm_interconnect_1_pio_key_s1_write_ports_inv <= not mm_interconnect_1_pio_key_s1_write;

	mm_interconnect_1_g_sensor_int_s1_write_ports_inv <= not mm_interconnect_1_g_sensor_int_s1_write;

	mm_interconnect_1_i2c_sda_s1_write_ports_inv <= not mm_interconnect_1_i2c_sda_s1_write;

	mm_interconnect_1_i2c_scl_s1_write_ports_inv <= not mm_interconnect_1_i2c_scl_s1_write;

	mm_interconnect_1_ext_sensor_int_s1_write_ports_inv <= not mm_interconnect_1_ext_sensor_int_s1_write;

	mm_interconnect_1_i2c_ext_sda_s1_write_ports_inv <= not mm_interconnect_1_i2c_ext_sda_s1_write;

	mm_interconnect_1_xbee_uart_s1_read_ports_inv <= not mm_interconnect_1_xbee_uart_s1_read;

	mm_interconnect_1_xbee_uart_s1_write_ports_inv <= not mm_interconnect_1_xbee_uart_s1_write;

	mm_interconnect_1_adc_spi_int_spi_control_port_read_ports_inv <= not mm_interconnect_1_adc_spi_int_spi_control_port_read;

	mm_interconnect_1_adc_spi_int_spi_control_port_write_ports_inv <= not mm_interconnect_1_adc_spi_int_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of DE0_nano_system
